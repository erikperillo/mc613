LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY demo_setup IS
	PORT (SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0) ;
		KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0) ;
		CLOCK_27: IN STD_LOGIC;
		CLOCK_50: IN STD_LOGIC;
		CLOCK_24: IN STD_LOGIC;
		EXT_CLOCK: IN STD_LOGIC;
		LEDR : OUT STD_LOGIC_VECTOR(0 TO 9) ;
		LEDG : OUT STD_LOGIC_VECTOR(0 TO 7) ;
		HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6) ;
		HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6) ;
		HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6) ;
		HEX3 : OUT STD_LOGIC_VECTOR(0 TO 6) );
END demo_setup ;

ARCHITECTURE Behavior OF demo_setup IS
BEGIN
	WITH SW SELECT
	HEX3 <= "0000001" WHEN "0000",
		"1001111" WHEN "0001",
		"0010010" WHEN "0010",
		"0000110" WHEN "0011",
		"1001100" WHEN "0100",
		"0100100" WHEN "0101",
		"0100000" WHEN "0110",
		"0001111" WHEN "0111",
		"0000000" WHEN "1000",
		"0000100" WHEN "1001",
		"0110000" WHEN OTHERS ;
END Behavior ;
